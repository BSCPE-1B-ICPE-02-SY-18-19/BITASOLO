CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 70 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 1477 636 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5283 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 971 252 0 3 22
0 4 5 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6874 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 649 243 0 3 22
0 16 15 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5305 0 0
2
5.89883e-315 0
0
2 +V
167 253 308 0 1 3
0 13
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
34 0 0
2
5.89883e-315 0
0
6 74LS48
188 1387 387 0 14 29
0 17 5 15 16 18 19 6 7 8
9 10 11 12 20
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
969 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 1387 670 0 17 19
10 12 11 10 9 8 7 6 21 2
0 1 1 0 0 0 0 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8402 0 0
2
5.89883e-315 0
0
6 74112~
219 1079 388 0 7 32
0 13 14 3 14 13 22 17
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3751 0 0
2
5.89883e-315 0
0
6 74112~
219 767 396 0 7 32
0 13 4 3 4 13 23 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
4292 0 0
2
5.89883e-315 0
0
6 74112~
219 523 397 0 7 32
0 13 16 3 16 13 24 15
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
6118 0 0
2
5.89883e-315 0
0
6 74112~
219 253 396 0 7 32
0 13 13 3 13 13 25 16
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
34 0 0
2
5.89883e-315 0
0
7 Pulser~
4 57 441 0 10 12
0 26 27 3 28 0 0 5 5 2
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6357 0 0
2
5.89883e-315 0
0
36
3 0 3 0 0 8192 0 8 0 0 36 3
737 369
629 369
629 514
9 1 2 0 0 8320 0 6 1 0 0 4
1387 628
1387 609
1477 609
1477 630
2 0 4 0 0 4096 0 8 0 0 4 2
743 360
670 360
3 4 4 0 0 4096 0 3 8 0 0 3
670 243
670 378
743 378
7 2 5 0 0 8192 0 8 2 0 0 4
791 360
871 360
871 261
947 261
7 7 6 0 0 8320 0 5 6 0 0 5
1419 351
1529 351
1529 765
1402 765
1402 706
8 6 7 0 0 8320 0 5 6 0 0 5
1419 360
1539 360
1539 755
1396 755
1396 706
9 5 8 0 0 8320 0 5 6 0 0 5
1419 369
1547 369
1547 747
1390 747
1390 706
10 4 9 0 0 8320 0 5 6 0 0 5
1419 378
1555 378
1555 736
1384 736
1384 706
11 3 10 0 0 8320 0 5 6 0 0 5
1419 387
1565 387
1565 729
1378 729
1378 706
12 2 11 0 0 8320 0 5 6 0 0 5
1419 396
1575 396
1575 719
1372 719
1372 706
13 1 12 0 0 8320 0 5 6 0 0 5
1419 405
1583 405
1583 711
1366 711
1366 706
0 0 13 0 0 4096 0 0 0 31 16 2
353 324
353 469
0 5 13 0 0 4224 0 0 7 15 0 3
767 469
1079 469
1079 400
0 5 13 0 0 0 0 0 8 16 0 3
523 469
767 469
767 408
5 5 13 0 0 0 0 10 9 0 0 4
253 408
253 469
523 469
523 409
2 0 14 0 0 4096 0 7 0 0 18 2
1055 352
1017 352
3 4 14 0 0 8320 0 2 7 0 0 4
992 252
1017 252
1017 370
1055 370
7 2 15 0 0 8192 0 9 3 0 0 4
547 361
594 361
594 252
625 252
0 7 16 0 0 8192 0 0 10 27 0 3
467 361
467 360
277 360
7 1 17 0 0 12416 0 7 5 0 0 5
1103 352
1103 593
1243 593
1243 351
1355 351
7 2 5 0 0 8320 0 8 5 0 0 5
791 360
791 611
1261 611
1261 360
1355 360
7 3 15 0 0 8320 0 9 5 0 0 5
547 361
547 631
1277 631
1277 369
1355 369
7 4 16 0 0 8320 0 10 5 0 0 5
277 360
277 647
1295 647
1295 378
1355 378
3 1 4 0 0 4224 0 3 2 0 0 2
670 243
947 243
3 0 3 0 0 0 0 9 0 0 36 3
493 370
423 370
423 514
2 0 16 0 0 0 0 9 0 0 28 2
499 361
467 361
4 1 16 0 0 0 0 9 3 0 0 4
499 379
467 379
467 234
625 234
1 0 13 0 0 0 0 7 0 0 30 2
1079 325
767 325
1 0 13 0 0 0 0 8 0 0 31 3
767 333
767 324
523 324
0 1 13 0 0 0 0 0 9 32 0 3
253 324
523 324
523 334
1 1 13 0 0 0 0 10 4 0 0 2
253 333
253 317
2 0 13 0 0 0 0 10 0 0 34 2
229 360
199 360
4 1 13 0 0 0 0 10 10 0 0 4
229 378
199 378
199 333
253 333
3 0 3 0 0 0 0 10 0 0 36 3
223 369
163 369
163 514
3 3 3 0 0 12416 0 11 7 0 0 6
81 432
115 432
115 514
990 514
990 361
1049 361
3
-35 0 0 0 400 255 0 0 0 3 2 1 34
15 Eras Medium ITC
0 0 0 30
507 144 1109 201
531 155 1084 196
30 BINARY 4 - BIT  SYNCHRONOUS UP
-35 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 23
150 17 607 81
176 29 580 73
23 Bitasolo, Shiela Mae L.
-29 0 0 0 400 255 0 0 0 3 2 1 18
8 Elephant
0 0 0 10
165 64 373 117
179 75 358 112
10 BSCpE - 1B
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
